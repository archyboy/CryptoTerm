module constants

pub const db_file_path = 'db/user.json'
