module constants

pub const db_file_path = 'src/db/user.json'
