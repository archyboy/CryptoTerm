module login
