module main

fn help_me(h string) {
	println('Help me with VLang please!!!')
}

fn thank_you(h string) {
	help_me('wææææ')
	println('Thanks you so much VLang :)')
}
