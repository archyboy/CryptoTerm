module config

pub struct Config {
pub mut:
	app_name    string = 'CryptoTerm'
	app_version string = '0.0.1'
}
