module main

fn help_me(msg string) {
	println(msg)
}

fn thank_you() {
	help_me('Thanks you so much VLang :)')
}
